/**
 * And gate: 
 * out = 1 if (a == 1 and b == 1)
 *       0 otherwise
 */

`default_nettype none
module And(
	input a,
	input b,
	output out
);
  wire w1;
  Nand NAND(.a(a), .b(b), .out(w1));
  Not NOT(.in(w1), .out(out));
endmodule
